// DE0_80MHZ.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module DE0_80MHZ (
		input  wire  ref_clk_clk,        //      ref_clk.clk
		input  wire  ref_reset_reset,    //    ref_reset.reset
		output wire  reset_source_reset, // reset_source.reset
		output wire  sys_clk_clk         //      sys_clk.clk
	);

	DE0_80MHZ_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (sys_clk_clk),        //      sys_clk.clk
		.reset_source_reset (reset_source_reset)  // reset_source.reset
	);

endmodule
